module not1(b,a);
output b;
input a;
assign b = ~a;
endmodule
